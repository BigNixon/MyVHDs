library ieee;
use ieee.std_logic_1164.all;

package ram_pkg is
    type memory is array(integer range <>) of std_logic_vector;
end package;

package body ram_pkg is
end package body;