library ieee;
use ieee.std_logic_1164.all;

package muxPackage is
    -- an array is a <n> group of std logic vector(any width)
    type mux_array is array (integer range <>) of std_logic_vector;

end muxPackage;


package body muxPackage is
end package body;